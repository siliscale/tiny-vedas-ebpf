typedef struct packed {
	logic alu;
	logic rs1;
	logic rs2;
	logic imm;
	logic rd;
	logic pc;
	logic load;
	logic store;
	logic lsu;
	logic add;
	logic sub;
	logic land;
	logic lor;
	logic lxor;
	logic sll;
	logic sra;
	logic srl;
	logic slt;
	logic unsign;
	logic condbr;
	logic beq;
	logic bne;
	logic bge;
	logic blt;
	logic bgt;
	logic jal;
	logic by;
	logic half;
	logic word;
	logic mul;
	logic rs1_sign;
	logic rs2_sign;
	logic low;
	logic divu;
	logic remu;
	logic nop;
	logic legal;
	logic offset;
	logic atomic;
	logic call;
	logic exit;
	logic arsh;
} decode_out_t;
